------------------------------------------------------------------
--Copyright 2017 Andrey S. Ionisyan (anserion@gmail.com)
--Licensed under the Apache License, Version 2.0 (the "License");
--you may not use this file except in compliance with the License.
--You may obtain a copy of the License at
--    http://www.apache.org/licenses/LICENSE-2.0
--Unless required by applicable law or agreed to in writing, software
--distributed under the License is distributed on an "AS IS" BASIS,
--WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--See the License for the specific language governing permissions and
--limitations under the License.
------------------------------------------------------------------

----------------------------------------------------------------------------------
-- Engineer: Andrey S. Ionisyan <anserion@gmail.com>
-- 
-- Description: vgafont ROM 8x16 patterns
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity rom_vgafont is
    Port ( 
		clk       : in STD_LOGIC;
		en        : in STD_LOGIC;
		addr      : in STD_LOGIC_VECTOR(11 downto 0);
		data      : out STD_LOGIC_VECTOR(7 downto 0)
	 );
end rom_vgafont;

architecture ax309 of rom_vgafont is
   type rom_type is array (0 to 4095) of std_logic_vector(7 downto 0);
   constant ROM : rom_type:= (
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"7E",x"81",x"A5",x"A5",x"A5",x"81",x"81",x"BD",x"99",x"81",x"7E",x"00",x"00",x"00",
x"00",x"00",x"7E",x"FF",x"DB",x"DB",x"DB",x"FF",x"FF",x"C3",x"E7",x"FF",x"7E",x"00",x"00",x"00",
x"00",x"00",x"6C",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"7C",x"38",x"10",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"10",x"38",x"7C",x"FE",x"7C",x"38",x"10",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"3C",x"3C",x"E7",x"E7",x"E7",x"18",x"18",x"3C",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"3C",x"7E",x"FF",x"FF",x"7E",x"18",x"18",x"3C",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"18",x"3C",x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E7",x"C3",x"C3",x"E7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"42",x"42",x"66",x"3C",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"C3",x"99",x"BD",x"BD",x"99",x"C3",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"1E",x"0E",x"1A",x"32",x"78",x"CC",x"CC",x"CC",x"78",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"3C",x"66",x"66",x"66",x"3C",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"3F",x"33",x"3F",x"30",x"30",x"30",x"70",x"F0",x"E0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"7F",x"63",x"7F",x"63",x"63",x"63",x"67",x"E7",x"E6",x"C0",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"18",x"DB",x"3C",x"E7",x"3C",x"DB",x"18",x"18",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"80",x"C0",x"E0",x"F8",x"FE",x"F8",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"02",x"06",x"0E",x"3E",x"FE",x"3E",x"0E",x"06",x"02",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"7E",x"3C",x"18",x"00",
x"00",x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"66",x"00",x"66",x"66",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"7F",x"DB",x"DB",x"DB",x"7B",x"1B",x"1B",x"1B",x"1B",x"00",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"60",x"38",x"6C",x"C6",x"C6",x"6C",x"38",x"0C",x"C6",x"7C",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"FE",x"FE",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"7E",x"3C",x"18",x"7E",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"7E",x"3C",x"18",x"00",
x"00",x"00",x"00",x"00",x"00",x"18",x"0C",x"FE",x"0C",x"18",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"30",x"60",x"FE",x"60",x"30",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"C0",x"C0",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"28",x"6C",x"FE",x"6C",x"28",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"10",x"38",x"38",x"7C",x"7C",x"FE",x"FE",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FE",x"7C",x"38",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"18",x"3C",x"3C",x"3C",x"3C",x"18",x"18",x"18",x"00",x"00",x"18",x"00",x"00",x"00",
x"00",x"66",x"66",x"66",x"66",x"66",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"6C",x"6C",x"6C",x"FE",x"6C",x"6C",x"6C",x"FE",x"6C",x"6C",x"6C",x"00",x"00",x"00",
x"18",x"18",x"18",x"7C",x"C6",x"C2",x"C0",x"7C",x"06",x"86",x"C6",x"7C",x"18",x"18",x"18",x"00",
x"00",x"00",x"00",x"00",x"00",x"C2",x"C6",x"0C",x"18",x"30",x"66",x"C6",x"00",x"00",x"00",x"00",
x"00",x"00",x"38",x"6C",x"6C",x"6C",x"38",x"76",x"DC",x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",
x"00",x"30",x"30",x"30",x"30",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"0C",x"18",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"18",x"0C",x"00",x"00",x"00",
x"00",x"00",x"30",x"18",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"18",x"30",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"66",x"66",x"3C",x"FF",x"3C",x"66",x"66",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"7E",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"30",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",
x"00",x"00",x"00",x"02",x"06",x"0C",x"18",x"30",x"60",x"C0",x"80",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"CE",x"DE",x"F6",x"F6",x"E6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"18",x"18",x"38",x"78",x"18",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"06",x"06",x"0C",x"18",x"30",x"60",x"C6",x"FE",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"06",x"06",x"06",x"3C",x"06",x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"0C",x"1C",x"3C",x"6C",x"CC",x"CC",x"FE",x"0C",x"0C",x"0C",x"1E",x"00",x"00",x"00",
x"00",x"00",x"FE",x"C0",x"C0",x"C0",x"FC",x"06",x"06",x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"38",x"60",x"C0",x"C0",x"FC",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"FE",x"C6",x"C6",x"06",x"06",x"0C",x"18",x"30",x"30",x"30",x"30",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"06",x"0C",x"78",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",
x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"30",x"00",x"00",
x"00",x"00",x"00",x"06",x"0C",x"18",x"30",x"60",x"30",x"18",x"0C",x"06",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"60",x"30",x"18",x"0C",x"06",x"0C",x"18",x"30",x"60",x"00",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"0C",x"18",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"DE",x"DE",x"DE",x"DC",x"C0",x"C0",x"7C",x"00",x"00",x"00",
x"00",x"00",x"10",x"38",x"6C",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"66",x"7C",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"C0",x"C0",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"FE",x"66",x"62",x"60",x"68",x"78",x"68",x"68",x"62",x"66",x"FE",x"00",x"00",x"00",
x"00",x"00",x"FE",x"66",x"62",x"60",x"68",x"78",x"68",x"68",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"C0",x"DE",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"3C",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"1E",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"CC",x"CC",x"78",x"00",x"00",x"00",
x"00",x"00",x"E6",x"66",x"66",x"6C",x"6C",x"78",x"6C",x"6C",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"F0",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"62",x"66",x"FE",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"E6",x"F6",x"FE",x"DE",x"CE",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"66",x"66",x"7C",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"D6",x"DE",x"7C",x"0C",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"66",x"7C",x"6C",x"66",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"60",x"38",x"0C",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"7E",x"7E",x"5A",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"6C",x"38",x"10",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"D6",x"D6",x"FE",x"7C",x"6C",x"6C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"6C",x"38",x"38",x"38",x"6C",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"3C",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"FE",x"C6",x"C6",x"8C",x"18",x"30",x"60",x"C2",x"C6",x"C6",x"FE",x"00",x"00",x"00",
x"00",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"80",x"C0",x"E0",x"70",x"38",x"1C",x"0E",x"06",x"02",x"00",x"00",x"00",x"00",
x"00",x"00",x"3C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"00",x"00",
x"10",x"10",x"38",x"6C",x"C6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",
x"30",x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"78",x"CC",x"0C",x"7C",x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",
x"00",x"00",x"E0",x"60",x"60",x"60",x"78",x"6C",x"66",x"66",x"66",x"66",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"1C",x"0C",x"0C",x"0C",x"3C",x"6C",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"FE",x"C0",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"38",x"6C",x"64",x"60",x"F0",x"60",x"60",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"76",x"CC",x"CC",x"CC",x"CC",x"CC",x"7C",x"0C",x"CC",x"78",x"00",
x"00",x"00",x"E0",x"60",x"60",x"6C",x"76",x"66",x"66",x"66",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"18",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"06",x"06",x"00",x"0E",x"06",x"06",x"06",x"06",x"06",x"06",x"66",x"66",x"3C",x"00",
x"00",x"00",x"E0",x"60",x"60",x"66",x"66",x"6C",x"78",x"6C",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"EC",x"FE",x"D6",x"D6",x"D6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"66",x"66",x"66",x"66",x"66",x"66",x"7C",x"60",x"F0",x"00",
x"00",x"00",x"00",x"00",x"00",x"76",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"7C",x"0C",x"1E",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"76",x"66",x"60",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"70",x"1C",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"10",x"30",x"30",x"FC",x"30",x"30",x"30",x"30",x"30",x"36",x"1C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"66",x"66",x"66",x"66",x"66",x"66",x"3C",x"18",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"D6",x"D6",x"FE",x"6C",x"6C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"6C",x"38",x"38",x"6C",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"0C",x"F8",x"00",
x"00",x"00",x"00",x"00",x"00",x"FE",x"C6",x"CC",x"18",x"30",x"66",x"C6",x"FE",x"00",x"00",x"00",
x"00",x"0E",x"18",x"18",x"18",x"18",x"18",x"70",x"70",x"18",x"18",x"18",x"18",x"18",x"0E",x"00",
x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"00",x"00",
x"00",x"70",x"18",x"18",x"18",x"18",x"18",x"0E",x"0E",x"18",x"18",x"18",x"18",x"18",x"70",x"00",
x"00",x"00",x"76",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"10",x"38",x"6C",x"C6",x"C6",x"C6",x"C6",x"FE",x"00",x"00",x"00",x"00",
x"00",x"00",x"10",x"38",x"6C",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"FE",x"66",x"62",x"60",x"7C",x"66",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"7C",x"66",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"FE",x"66",x"62",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"3E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"FF",x"C3",x"C3",x"00",
x"00",x"00",x"FE",x"66",x"66",x"62",x"68",x"78",x"68",x"62",x"66",x"66",x"FE",x"00",x"00",x"00",
x"00",x"00",x"D6",x"D6",x"D6",x"7C",x"38",x"7C",x"D6",x"D6",x"D6",x"D6",x"D6",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"06",x"06",x"06",x"3C",x"06",x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"CE",x"DE",x"FE",x"F6",x"E6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"38",x"38",x"C6",x"C6",x"CE",x"DE",x"FE",x"F6",x"E6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"E6",x"66",x"6C",x"6C",x"78",x"6C",x"6C",x"66",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"3E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"FE",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"FC",x"66",x"66",x"66",x"66",x"66",x"7C",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"C0",x"C0",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"7E",x"7E",x"5A",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"06",x"06",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"18",x"7E",x"DB",x"DB",x"DB",x"DB",x"DB",x"DB",x"DB",x"7E",x"18",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"6C",x"38",x"38",x"38",x"6C",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FE",x"06",x"06",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"06",x"06",x"06",x"00",x"00",x"00",
x"00",x"00",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"FE",x"00",x"00",x"00",
x"00",x"00",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"FE",x"03",x"03",x"00",
x"00",x"00",x"F8",x"F0",x"B0",x"30",x"3C",x"36",x"36",x"36",x"36",x"36",x"7C",x"00",x"00",x"00",
x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"F6",x"DE",x"DE",x"DE",x"DE",x"DE",x"F6",x"00",x"00",x"00",
x"00",x"00",x"F0",x"60",x"60",x"60",x"7C",x"66",x"66",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"78",x"CC",x"86",x"86",x"26",x"3E",x"26",x"86",x"86",x"CC",x"78",x"00",x"00",x"00",
x"00",x"00",x"9C",x"B6",x"B6",x"B6",x"B6",x"F6",x"B6",x"B6",x"B6",x"B6",x"9C",x"00",x"00",x"00",
x"00",x"00",x"7E",x"CC",x"CC",x"CC",x"CC",x"7C",x"6C",x"CC",x"CC",x"CE",x"CE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"78",x"CC",x"0C",x"7C",x"CC",x"CC",x"CC",x"76",x"00",x"00",x"00",
x"00",x"00",x"00",x"1C",x"30",x"60",x"7C",x"66",x"66",x"66",x"66",x"66",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FC",x"66",x"66",x"7C",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FE",x"62",x"60",x"60",x"60",x"60",x"60",x"F0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"3E",x"66",x"66",x"66",x"66",x"66",x"66",x"FF",x"C3",x"C3",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"FE",x"C0",x"C0",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"7C",x"7C",x"D6",x"D6",x"D6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"66",x"0C",x"06",x"66",x"66",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"CE",x"DE",x"FE",x"F6",x"E6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"38",x"38",x"00",x"C6",x"CE",x"DE",x"FE",x"F6",x"E6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E6",x"66",x"6C",x"78",x"6C",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"3E",x"66",x"66",x"66",x"66",x"66",x"66",x"E6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"EE",x"FE",x"FE",x"D6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"FE",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FE",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"00",x"00",x"00",
x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",x"44",x"11",
x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",
x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",x"77",x"DD",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"F6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"18",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"36",x"36",x"36",x"36",x"36",x"36",x"F6",x"06",x"F6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"06",x"F6",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"F6",x"06",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"18",x"18",x"18",x"18",x"18",x"18",x"F8",x"18",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"30",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"F7",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"F7",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"37",x"30",x"37",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"36",x"36",x"36",x"36",x"36",x"36",x"F7",x"00",x"F7",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"3F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"18",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"18",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3F",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"36",x"FF",x"36",x"36",x"36",x"36",x"36",x"36",x"36",
x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"18",x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"DC",x"66",x"66",x"66",x"66",x"66",x"7C",x"60",x"60",x"F0",x"00",
x"00",x"00",x"00",x"00",x"00",x"7C",x"C6",x"C6",x"C0",x"C0",x"C6",x"C6",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7E",x"5A",x"18",x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"0C",x"F8",x"00",
x"00",x"00",x"00",x"00",x"00",x"18",x"7E",x"DB",x"DB",x"DB",x"DB",x"DB",x"7E",x"18",x"18",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"6C",x"38",x"38",x"6C",x"C6",x"C6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FE",x"06",x"06",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"C6",x"C6",x"7E",x"06",x"06",x"06",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"FE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"D6",x"FE",x"03",x"03",x"00",
x"00",x"00",x"00",x"00",x"00",x"F8",x"B0",x"3C",x"36",x"36",x"36",x"36",x"7C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"C6",x"C6",x"F6",x"DE",x"DE",x"DE",x"DE",x"F6",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"F0",x"60",x"60",x"7C",x"66",x"66",x"66",x"FC",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"06",x"1E",x"06",x"66",x"66",x"3C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"9C",x"B6",x"B6",x"F6",x"B6",x"B6",x"B6",x"9C",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"7E",x"CC",x"CC",x"CC",x"7C",x"6C",x"CC",x"CE",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"FE",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"30",x"18",x"0C",x"06",x"0C",x"18",x"30",x"00",x"7E",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"0C",x"18",x"30",x"60",x"30",x"18",x"0C",x"00",x"7E",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"0E",x"1B",x"1B",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"D8",x"D8",x"70",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"7E",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"76",x"DC",x"00",x"76",x"DC",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"38",x"6C",x"6C",x"6C",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"0F",x"0C",x"0C",x"0C",x"0C",x"0C",x"EC",x"6C",x"3C",x"1C",x"0C",x"00",x"00",x"00",x"00",
x"00",x"00",x"D8",x"6C",x"6C",x"6C",x"6C",x"6C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"70",x"D8",x"30",x"60",x"C8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
);
   signal rdata: std_logic_vector(7 downto 0);
begin
	rdata<=ROM(conv_integer(addr));
   process(clk)
   begin
		if rising_edge(clk) then
         if en='1' then
            data<=rdata;
         end if;
		end if;
	end process;
end ax309;